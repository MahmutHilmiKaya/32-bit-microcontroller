library IEEE;
use IEEE.STD_LOGIC_1164.ALL;


////////////////////////////////////////////////////////////////////////////////
// Last Edits: Dr. Burak Unal
// 
// Module - PCAdder.vhd
// Description - 32-Bit program counter (PC) adder.
// 
// INPUTS:-
// PCResult: 32-Bit input port.
// 
// OUTPUTS:-
// PCAddResult: 32-Bit output port.
//
// FUNCTIONALITY:-
// Design an incrementor by 4 
// (a hard-wired ADDER whose first input is from the PCResult, and 
// whose second input is a hard-wired value of 4 that outputs PCResult + 4. 
// The result should always be an increment of the signal 'PCResult' by 4 (i.e., PCAddResult = PCResult + 4).
////////////////////////////////////////////////////////////////////////////////


